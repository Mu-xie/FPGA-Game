----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    13:41:17 05/12/2015 
-- Design Name: 
-- Module Name:    obstacles2_ROM - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity obstacles2_ROM is
    Port ( obstacle2_on     : in  STD_LOGIC;
           obstacle2_row    : in  STD_LOGIC_VECTOR (10 downto 0);
           obstacle2_col    : in  STD_LOGIC_VECTOR (9 downto 0);
			  obstacle2_enable : out  STD_LOGIC;
           obstacle2_rgb    : out  STD_LOGIC );
end obstacles2_ROM;

architecture Behavioral of obstacles2_ROM is
type ROM is array(0 to 49) of std_logic_vector(49 downto 0);
constant content : ROM := (
 0 => "00000000000000000000000000000000000000000000000000",
 1 => "00000000000000000000000000000000000000000000000000",
 2 => "00000000000000000000000000000000000000000000000000",
 3 => "00000000000000000000000000000000000000000000000000",
 4 => "00000000000000000000000000000000000000000000000000",
 5 => "00000000000000000000000000011000000000000000000000",
 6 => "00000000000000000000000000011110000000000000000000",
 7 => "00000000000000000100000001111111100000000000000000",
 8 => "00000000000000011110000011111111110000000000000000",
 9 => "00000000000001111111011111111111111111000000000000",
10 => "00000000000011111111111111111111111111110000000000",
11 => "00000000001111111111111111111111111111111100000000",
12 => "00000001111111111111111111111111111111111000000000",
13 => "00000001111111111111111111111111111111110000000000",
14 => "00000001111111111111111111111111111111110000000000",
15 => "00000000111111111111111111111111111111111110000000",
16 => "00000000111111111111111111111111111111111111111000",
17 => "00000000011111111111111111111111111111111111111000",
18 => "00000000111111111111111111111111111111111111111100",
19 => "00000000111111111111111111111111111110001111111100",
20 => "00000001111111111101111111111111111100000111111110",
21 => "00000011111111111000111111111111111100000111111110",
22 => "00000111111111111000011111111111111110001111111100",
23 => "00000011111111111100111111111111111111111111111000",
24 => "00000001111111111111111111111111111111111111110000",
25 => "00000000111111111111111111111111111111111111100000",
26 => "00000000111111111111111111111111111111111110000000",
27 => "00000000011111111111111111111111111111111110000000",
28 => "00000000001111111111111111111111111111111100000000",
29 => "00000000111111111111111111111111111111111100000000",
30 => "00000000111111111111111111111111111111111000000000",
31 => "00000000001111111111111111111111111111110000000000",
32 => "00000000001111111111111111111111111110000000000000",
33 => "00000000000111111111111111111111111110000000000000",
34 => "00000000001111111111000000011110000000000000000000",
35 => "00000000000001111000000000000000000000000000000000",
36 => "00000000000000000000000000000000000000000000000000",
37 => "00000000000000000000000000000000000000000000000000",
38 => "00000000000000000000000000000000000000000000000000",
39 => "00000000000000000000000000000000000000000000000000",
40 => "00000000000000000000000000000000000000000000000000",
41 => "00000000000000000000000000000000000000000000000000",
42 => "00000000000000000000000000000000000000000000000000",
43 => "00000000000000000000000000000000000000000000000000",
44 => "00000000000000000000000000000000000000000000000000",
45 => "00000000000000000000000000000000000000000000000000",
46 => "00000000000000000000000000000000000000000000000000",
47 => "00000000000000000000000000000000000000000000000000",
48 => "00000000000000000000000000000000000000000000000000",
49 => "00000000000000000000000000000000000000000000000000"
	);

signal data_line : std_logic_vector(0 to 49);
signal obs2_rgb : std_logic;
signal enable : std_logic;
constant rest : integer := 2;
begin

process(obstacle2_on, obstacle2_col, data_line, obstacle2_row)
begin

    obs2_rgb <= '0';
	 enable <= '0';
	 
    -- IF OBSTACLE IS ON
    if obstacle2_on = '1' then
	     -- SCALING ALGORITHM
		  if (conv_integer(obstacle2_col) rem rest) = 0 then
	         data_line <= content((conv_integer(obstacle2_col)) / rest);
		  else
		      data_line <= content((conv_integer(obstacle2_col) - (conv_integer(obstacle2_col) rem rest)) / rest);
		  end if;
		  if (conv_integer(obstacle2_row) rem rest) = 0 then
		      obs2_rgb <= data_line((conv_integer(obstacle2_row)) / rest);
				-- ENABLE ROM
				enable <= '1';
		  else
		  		obs2_rgb <= data_line((conv_integer(obstacle2_row) - (conv_integer(obstacle2_row) rem rest)) / rest);
				-- ENABLE ROM
				enable <= '1';
		  end if;
	 end if;

end process;

obstacle2_rgb <= obs2_rgb;
obstacle2_enable <= enable;

end Behavioral;