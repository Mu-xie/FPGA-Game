----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    11:44:13 05/21/2015 
-- Design Name: 
-- Module Name:    shoot_ROM - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity shoot_ROM is
    Port ( shoot_on  : in  STD_LOGIC;
           shoot_row : in  STD_LOGIC_VECTOR (10 downto 0);
           shoot_col : in  STD_LOGIC_VECTOR (9 downto 0);
           shoot_rgb : out  STD_LOGIC );
end shoot_ROM;

architecture Behavioral of shoot_ROM is
type ROM is array(0 to 39) of std_logic_vector(39 downto 0);
constant content : ROM := (
 0 => "0000000000000000000110000000000000000000",
 1 => "0000000000000000001111000000000000000000",
 2 => "0011110000000000011001100000000000111100",
 3 => "0010001100000000110000110000000011000100",
 4 => "0010000010000000110000110000000100000100",
 5 => "0010011111111111111111111111111111100100",
 6 => "0001010001111111111111111111111000101000",
 7 => "0001010011000000000000000000001100101000",
 8 => "0000110110000000000000000000000110110000",
 9 => "0000011100111111111111111111110011100000",
10 => "0000011001111111111111111111111001100000",
11 => "0000011001111111111111111111111001100000",
12 => "0000011001111111111111111111111001100000",
13 => "0000011001111111111111111111111001100000",
14 => "0000011001111111111111111111111001100000",
15 => "0000011001111111111111111111111001100000",
16 => "0001111001111111111111111111111001111000",
17 => "0011111001111111111001111111111001111100",
18 => "0110011001111111110000111111111001100110",
19 => "1100011001111111100000011111111001100011",
20 => "1100011001111111100000011111111001100011",
21 => "0110011001111111110000111111111001100110",
22 => "0011111001111111111001111111111001111100",
23 => "0001111001111111111111111111111001111000",
24 => "0000011001111111111111111111111001100000",
25 => "0000011001111111111111111111111001100000",
26 => "0000011001111111111111111111111001100000",
27 => "0000011001111111111111111111111001100000",
28 => "0000011001111111111111111111111001100000",
29 => "0000011001111111111111111111111001100000",
30 => "0000011100111111111111111111110011100000",
31 => "0000110110000000000000000000000110110000",
32 => "0001010011000000000000000000001100101000",
33 => "0001010001111111111111111111111000101000",
34 => "0010011111111111111111111111111111100100",
35 => "0010000010000000110000110000000100000100",
36 => "0010001100000000110000110000000011000100",
37 => "0011110000000000011001100000000000111100",
38 => "0000000000000000001111000000000000000000",
39 => "0000000000000000000110000000000000000000"
);
signal data_line : std_logic_vector(0 to 39);
signal rgb : std_logic;
begin

process(shoot_on, shoot_col, data_line, shoot_row)
begin

    rgb <= '0';

    if shoot_on = '1' then
		  	 data_line <= content(conv_integer(shoot_col));
	       rgb <= data_line(conv_integer(shoot_row));
	 end if;
	 
end process;

shoot_rgb <= rgb;

end Behavioral;









