----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    13:40:58 05/12/2015 
-- Design Name: 
-- Module Name:    obstacles1_ROM - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity obstacles1_ROM is
    Port ( obstacle1_on     : in  STD_LOGIC;
           obstacle1_row    : in  STD_LOGIC_VECTOR (10 downto 0);
           obstacle1_col    : in  STD_LOGIC_VECTOR (9 downto 0);
			  obstacle1_enable : out  STD_LOGIC;
           obstacle1_rgb    : out  STD_LOGIC );
end obstacles1_ROM;

architecture Behavioral of obstacles1_ROM is
type ROM is array(0 to 49) of std_logic_vector(49 downto 0);
constant content : ROM := (
 0 => "00000000000000000000000000000000000000000000000000",
 1 => "00000000000000000000000000000000000000000000000000",
 2 => "00000000000000000000000000000000000000000000000000",
 3 => "00000000000000000000000000000000000000000000000000",
 4 => "00000000000000000000000000000000000000000000000000",
 5 => "00000000000000000000000000000000000000111000000000",
 6 => "00000000000000000000000000000000000001111111100000",
 7 => "00000000000000000000000010000000000001111111111100",
 8 => "00000000000000000000011110001111001111111111111100",
 9 => "00000000000000000001111111011111111111111111111000",
10 => "00000000000000001111111111111111111111111111111000",
11 => "00000000000000111111111111111111111111111111111000",
12 => "00000000001111111111111111111111111111111111110000",
13 => "00000000001111111111111111111111111111111111110000",
14 => "00000000000111111111111111111111111111111111100000",
15 => "00000000000011111111111111111111111111111111100000",
16 => "00000000000011111111111100001111111111111111100000",
17 => "00000000000111111111111110001111111111111111100000",
18 => "00000000000111111111111110000111111111111111000000",
19 => "00000000001111111111111100001111111111111111000000",
20 => "00000000001111111111111111000111111111111111000000",
21 => "00000000001111111111111111111111111111111111100000",
22 => "00000000011111111111111111111111111111111111110000",
23 => "00000000111111111111111111111111111111111111111000",
24 => "00000001111111111111111111111111111111111111111100",
25 => "00000011111111111111111111111111111111001111111100",
26 => "00000111111111111111111111111111111110001011111100",
27 => "00000001111111111011111111111111111111000011111000",
28 => "00000001111111100000111111111111111111101111111000",
29 => "00000000111111000000011111111111111111111111111000",
30 => "00000000111111100000111111111111111111111100000000",
31 => "00000000111111111011111111111111111111111100000000",
32 => "00000000011111111111111111111110111111111100000000",
33 => "00000000000111111111111111110000011111110000000000",
34 => "00000000000001111111111110000000001111000000000000",
35 => "00000000000000011111110000000000000110000000000000",
36 => "00000000000000001111100000000000000000000000000000",
37 => "00000000000000000111000000000000000000000000000000",
38 => "00000000000000000010000000000000000000000000000000",
39 => "00000000000000000000000000000000000000000000000000",
40 => "00000000000000000000000000000000000000000000000000",
41 => "00000000000000000000000000000000000000000000000000",
42 => "00000000000000000000000000000000000000000000000000",
43 => "00000000000000000000000000000000000000000000000000",
44 => "00000000000000000000000000000000000000000000000000",
45 => "00000000000000000000000000000000000000000000000000",
46 => "00000000000000000000000000000000000000000000000000",
47 => "00000000000000000000000000000000000000000000000000",
48 => "00000000000000000000000000000000000000000000000000",
49 => "00000000000000000000000000000000000000000000000000"
	);

signal data_line : std_logic_vector(0 to 49);
signal obs1_rgb : std_logic;
signal enable : std_logic;
constant rest : integer := 2;
begin

process(obstacle1_on, obstacle1_col, obstacle1_row)
begin

    obs1_rgb <= '0';
	 enable <= '0';
	 
    -- IF OBSTACLE IS ON
    if obstacle1_on = '1' then
	     -- SCALING ALGORITHM
		  if (conv_integer(obstacle1_col) rem rest) = 0 then
	         data_line <= content((conv_integer(obstacle1_col)) / rest);
		  else
		      data_line <= content((conv_integer(obstacle1_col) - (conv_integer(obstacle1_col) rem rest)) / rest);
		  end if;
		  if (conv_integer(obstacle1_row) rem rest) = 0 then
		      obs1_rgb <= data_line((conv_integer(obstacle1_row)) / rest);
			   -- ENABLE ROM
				enable <= '1';
		  else
		  		obs1_rgb <= data_line((conv_integer(obstacle1_row) - (conv_integer(obstacle1_row) rem rest)) / rest);
				-- ENABLE ROM
				enable <= '1';
		  end if;
	 end if;

end process;

obstacle1_rgb <= obs1_rgb;
obstacle1_enable <= enable;

end Behavioral;